library ieee ;
use ieee.std_logic_1164.all;

package components is

  component CC_PLL
  generic (
    REF_CLK         : string := "0";          -- reference clk in MHz
    OUT_CLK         : string := "0";          -- output clk in MHz
    PERF_MD         : string := "UNDEFINED";  -- LOWPOWER, ECONOMY, SPEED (optional, global, setting of Place&Route can be used instead)
    LOW_JITTER      : natural := 1;           -- 0: disable, 1: enable low jitter mode
    CI_FILTER_CONST : natural := 2;           -- optional CI filter constant
    CP_FILTER_CONST : natural := 4            -- optional CP filter constant
  );
  port (
    CLK_REF             : in std_logic;
    CLK_FEEDBACK        : in std_logic;
    USR_CLK_REF         : in std_logic;
    USR_LOCKED_STDY_RST : in std_logic;
    USR_PLL_LOCKED_STDY : out std_logic;
    USR_PLL_LOCKED      : out std_logic;
    CLK270              : out std_logic;
    CLK180              : out std_logic;
    CLK0                : out std_logic;
    CLK90               : out std_logic;
    CLK_REF_OUT         : out std_logic
  );
  end component;

  component CC_PLL_ADV
  generic (
    PLL_CFG_A : std_logic_vector(95 downto 0) := (others => 'X');
    PLL_CFG_B : std_logic_vector(95 downto 0) := (others => 'X')
  );
  port (
    CLK_REF             : in std_logic;
    CLK_FEEDBACK        : in std_logic;
    USR_CLK_REF         : in std_logic;
    USR_LOCKED_STDY_RST : in std_logic;
    USR_SEL_A_B         : in std_logic;
    USR_PLL_LOCKED_STDY : out std_logic;
    USR_PLL_LOCKED      : out std_logic;
    CLK270              : out std_logic;
    CLK180              : out std_logic;
    CLK0                : out std_logic;
    CLK90               : out std_logic;
    CLK_REF_OUT         : out std_logic
  );
  end component;

  component CC_SERDES
  generic (
    SERDES_CFG : string := ""
  );
  port (
    TX_DATA_I             : in std_logic_vector(63 downto 0);
    TX_RESET_I            : in std_logic;
    TX_PCS_RESET_I        : in std_logic;
    TX_PMA_RESET_I        : in std_logic;
    PLL_RESET_I           : in std_logic;
    TX_POWERDOWN_N_I      : in std_logic;
    TX_POLARITY_I         : in std_logic;
    TX_PRBS_SEL_I         : in std_logic_vector(2 downto 0);
    TX_PRBS_FORCE_ERR_I   : in std_logic;
    TX_8B10B_EN_I         : in std_logic;
    TX_8B10B_BYPASS_I     : in std_logic_vector(7 downto 0);
    TX_CHAR_IS_K_I        : in std_logic_vector(7 downto 0);
    TX_CHAR_DISPMODE_I    : in std_logic_vector(7 downto 0);
    TX_CHAR_DISPVAL_I     : in std_logic_vector(7 downto 0);
    TX_ELEC_IDLE_I        : in std_logic;
    TX_DETECT_RX_I        : in std_logic;
    LOOPBACK_I            : in std_logic_vector(2 downto 0);
    CLK_CORE_TX_I         : in std_logic;
    CLK_CORE_RX_I         : in std_logic;
    RX_RESET_I            : in std_logic;
    RX_PMA_RESET_I        : in std_logic;
    RX_EQA_RESET_I        : in std_logic;
    RX_CDR_RESET_I        : in std_logic;
    RX_PCS_RESET_I        : in std_logic;
    RX_BUF_RESET_I        : in std_logic;
    RX_POWERDOWN_N_I      : in std_logic;
    RX_POLARITY_I         : in std_logic;
    RX_PRBS_SEL_I         : in std_logic_vector(2 downto 0);
    RX_PRBS_CNT_RESET_I   : in std_logic;
    RX_8B10B_EN_I         : in std_logic;
    RX_8B10B_BYPASS_I     : in std_logic_vector(7 downto 0);
    RX_EN_EI_DETECTOR_I   : in std_logic;
    RX_COMMA_DETECT_EN_I  : in std_logic;
    RX_SLIDE_I            : in std_logic;
    RX_MCOMMA_ALIGN_I     : in std_logic;
    RX_PCOMMA_ALIGN_I     : in std_logic;
    CLK_REG_I             : in std_logic;
    REGFILE_WE_I          : in std_logic;
    REGFILE_EN_I          : in std_logic;
    REGFILE_ADDR_I        : in std_logic_vector(7 downto 0);
    REGFILE_DI_I          : in std_logic_vector(15 downto 0);
    REGFILE_MASK_I        : in std_logic_vector(15 downto 0);
    RX_DATA_O            : out std_logic_vector(63 downto 0);
    RX_NOT_IN_TABLE_O    : out std_logic_vector(7 downto 0);
    RX_CHAR_IS_COMMA_O   : out std_logic_vector(7 downto 0);
    RX_CHAR_IS_K_O       : out std_logic_vector(7 downto 0);
    RX_DISP_ERR_O        : out std_logic_vector(7 downto 0);
    RX_DETECT_DONE_O     : out std_logic;
    RX_PRESENT_O         : out std_logic;
    TX_BUF_ERR_O         : out std_logic;
    TX_RESETDONE_O       : out std_logic;
    RX_PRBS_ERR_O        : out std_logic;
    RX_BUF_ERR_O         : out std_logic;
    RX_BYTE_IS_ALIGNED_O : out std_logic;
    RX_BYTE_REALIGN_O    : out std_logic;
    RX_RESETDONE_O       : out std_logic;
    RX_EI_EN_O           : out std_logic;
    CLK_CORE_RX_O        : out std_logic;
    CLK_CORE_PLL_O       : out std_logic;
    REGFILE_DO_O         : out std_logic_vector(15 downto 0);
    REGFILE_RDY_O        : out std_logic
  );
  end component;

  component CC_CFG_CTRL
  port (
    DATA  : in std_logic_vector(7 downto 0);
    CLK   : in std_logic;
    EN    : in std_logic;
    RECFG : in std_logic;
    VALID : in std_logic
  );
  end component;

  component CC_BRAM_20K is
  generic (
    -- Location format: D(0..N-1)X(0..3)Y(0..7) or UNPLACED
    LOC : string := "UNPLACED";
    -- Port Widths
    A_RD_WIDTH : natural := 0;
    B_RD_WIDTH : natural := 0;
    A_WR_WIDTH : natural := 0;
    B_WR_WIDTH : natural := 0;
    -- RAM and Write Modes
    RAM_MODE  : string := "SDP";
    A_WR_MODE : string := "NO_CHANGE";
    B_WR_MODE : string := "NO_CHANGE";
    -- Inverting Control Pins
    A_CLK_INV : std_logic := '0';
    B_CLK_INV : std_logic := '0';
    A_EN_INV  : std_logic := '0';
    B_EN_INV  : std_logic := '0';
    A_WE_INV  : std_logic := '0';
    B_WE_INV  : std_logic := '0';
    -- Output Register
    A_DO_REG : std_logic := '0';
    B_DO_REG : std_logic := '0';
    -- Error Checking and Correction
    ECC_EN : std_logic := '0';
    -- RAM init content
    INIT_00 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_01 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_02 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_03 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_04 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_05 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_06 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_07 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_08 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_09 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_10 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_11 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_12 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_13 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_14 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_15 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_16 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_17 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_18 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_19 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_20 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_21 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_22 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_23 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_24 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_25 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_26 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_27 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_28 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_29 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_30 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_31 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_32 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_33 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_34 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_35 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_36 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_37 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_38 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_39 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000"
  );
  port (
    -- clocks
    A_CLK        : in std_logic;
    B_CLK        : in std_logic;
    -- inputs
    A_EN         : in std_logic;
    B_EN         : in std_logic;
    A_WE         : in std_logic;
    B_WE         : in std_logic;
    A_ADDR       : in std_logic_vector(15 downto 0);
    B_ADDR       : in std_logic_vector(15 downto 0);
    A_DI         : in std_logic_vector(19 downto 0);
    B_DI         : in std_logic_vector(19 downto 0);
    A_BM         : in std_logic_vector(19 downto 0);
    B_BM         : in std_logic_vector(19 downto 0);
    -- outputs
    A_DO         : out std_logic_vector(19 downto 0);
    B_DO         : out std_logic_vector(19 downto 0);
    ECC_1B_ERR   : out std_logic;
    ECC_2B_ERR   : out std_logic
  );
  end component;

  component CC_BRAM_40K is
  generic (
    -- Location format: D(0..N-1)X(0..3)Y(0..7) or UNPLACED
    LOC : string := "UNPLACED";
    CAS : string := "NONE";      -- NONE, UPPER, LOWER
    -- Port Widths
    A_RD_WIDTH : natural := 0;
    B_RD_WIDTH : natural := 0;
    A_WR_WIDTH : natural := 0;
    B_WR_WIDTH : natural := 0;
    -- RAM and Write Modes
    RAM_MODE  : string := "SDP";
    A_WR_MODE : string := "NO_CHANGE";
    B_WR_MODE : string := "NO_CHANGE";
    -- Inverting Control Pins
    A_CLK_INV : std_logic := '0';
    B_CLK_INV : std_logic := '0';
    A_EN_INV  : std_logic := '0';
    B_EN_INV  : std_logic := '0';
    A_WE_INV  : std_logic := '0';
    B_WE_INV  : std_logic := '0';
    -- Output Register
    A_DO_REG : std_logic := '0';
    B_DO_REG : std_logic := '0';
    -- Error Checking and Correction
    A_ECC_EN : std_logic := '0';
    B_ECC_EN : std_logic := '0';
    -- RAM init content
    INIT_00 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_01 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_02 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_03 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_04 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_05 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_06 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_07 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_08 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_09 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_0F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_10 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_11 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_12 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_13 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_14 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_15 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_16 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_17 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_18 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_19 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_1F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_20 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_21 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_22 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_23 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_24 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_25 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_26 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_27 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_28 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_29 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_2F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_30 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_31 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_32 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_33 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_34 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_35 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_36 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_37 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_38 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_39 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_3F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_40 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_41 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_42 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_43 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_44 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_45 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_46 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_47 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_48 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_49 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_4A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_4B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_4C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_4D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_4E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_4F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_50 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_51 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_52 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_53 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_54 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_55 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_56 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_57 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_58 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_59 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_5A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_5B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_5C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_5D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_5E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_5F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_60 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_61 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_62 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_63 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_64 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_65 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_66 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_67 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_68 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_69 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_6A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_6B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_6C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_6D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_6E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_6F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_70 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_71 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_72 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_73 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_74 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_75 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_76 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_77 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_78 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_79 : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_7A : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_7B : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_7C : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_7D : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_7E : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    INIT_7F : std_logic_vector(319 downto 0) := x"00000000000000000000000000000000000000000000000000000000000000000000000000000000"
  );
  port (
    -- clocks
    A_CLK        : in std_logic;
    B_CLK        : in std_logic;
    -- inputs
    A_EN         : in std_logic;
    B_EN         : in std_logic;
    A_WE         : in std_logic;
    B_WE         : in std_logic;
    A_ADDR       : in std_logic_vector(15 downto 0);
    B_ADDR       : in std_logic_vector(15 downto 0);
    A_DI         : in std_logic_vector(39 downto 0);
    B_DI         : in std_logic_vector(39 downto 0);
    A_BM         : in std_logic_vector(39 downto 0);
    B_BM         : in std_logic_vector(39 downto 0);
    A_CI         : in std_logic;
    B_CI         : in std_logic;
    -- outputs
    A_DO         : out std_logic_vector(39 downto 0);
    B_DO         : out std_logic_vector(39 downto 0);
    A_ECC_1B_ERR : out std_logic;
    B_ECC_1B_ERR : out std_logic;
    A_ECC_2B_ERR : out std_logic;
    B_ECC_2B_ERR : out std_logic
    -- These ports are listed in the Primitives Doc, but p_r tool doesn't knows them:
    --   FATAL ERROR: (51513): Component CC_BRAM_40K has no port name: A_CO
    --   FATAL ERROR: (51513): Component CC_BRAM_40K has no port name: B_CO
--    A_CO         : out std_logic;
--    B_CO         : out std_logic
  );
  end component;

  component CC_FIFO_40K
    generic (
    LOC                 : string := "UNPLACED";  -- Location format: D(0..N-1)X(0..3)Y(0..7) or UNPLACED
    ALMOST_FULL_OFFSET  : std_logic_vector (12 downto 0) := (others => '0');  -- Almost full offset
    ALMOST_EMPTY_OFFSET : std_logic_vector (12 downto 0) := (others => '0');  -- Almost empty offset
    A_WIDTH             : natural := 0;      -- Port A Width
    B_WIDTH             : natural := 0;      -- Port B Width
    RAM_MODE            : string := "SDP";   -- RAM mode: "TPD" or "SDP"
    FIFO_MODE           : string := "SYNC";  -- Write mode: "ASYNC" or "SYNC"
    A_CLK_INV           : std_logic := '0';  -- Inverting Control Pins
    B_CLK_INV           : std_logic := '0';  -- Inverting Control Pins
    A_EN_INV            : std_logic := '0';  -- Inverting Control Pins
    B_EN_INV            : std_logic := '0';  -- Inverting Control Pins
    A_WE_INV            : std_logic := '0';  -- Inverting Control Pins
    B_WE_INV            : std_logic := '0';  -- Inverting Control Pins
    A_DO_REG            : std_logic := '0';  -- Port A Output Register
    B_DO_REG            : std_logic := '0';  -- Port B Output Register
    A_ECC_EN            : std_logic := '0';  -- Port A Error Checking and Correction
    B_ECC_EN            : std_logic := '0'   -- Port B Error Checking and Correction
    );
  port (
    A_ECC_1B_ERR : out std_logic;
    B_ECC_1B_ERR : out std_logic;
    A_ECC_2B_ERR : out std_logic;
    B_ECC_2B_ERR : out std_logic;
    -- FIFO pop port
    A_DO : out std_logic_vector(39 downto 0);
    B_DO : out std_logic_vector(39 downto 0);
  
    A_CLK : in std_logic;
    A_EN  : in std_logic;
    -- FIFO push port
    A_DI : in std_logic_vector(39 downto 0);
    B_DI : in std_logic_vector(39 downto 0);
    A_BM : in std_logic_vector(39 downto 0);
    B_BM : in std_logic_vector(39 downto 0);
  
    B_CLK : in std_logic;
    B_EN  : in std_logic;
    B_WE  : in std_logic;
    -- FIFO control
    F_RST_N : in std_logic;
    F_ALMOST_FULL_OFFSET  : in std_logic_vector(12 downto 0);
    F_ALMOST_EMPTY_OFFSET : in std_logic_vector(12 downto 0);
    -- FIFO status signals
    F_FULL         : out std_logic;
    F_EMPTY        : out std_logic;
    F_ALMOST_FULL  : out std_logic;
    F_ALMOST_EMPTY : out std_logic;
    F_RD_ERROR     : out std_logic;
    F_WR_ERROR     : out std_logic;
    F_RD_PTR       : out std_logic_vector(15 downto 0);
    F_WR_PTR       : out std_logic_vector(15 downto 0)
  );
  end component;

  component CC_CFG_END
  port (
    CFG_END : out std_logic
  );
  end component;

  component CC_BUFG
  port (
    I : in  std_logic;
    O : out std_logic
  );
  end component;


end package components;